module and_gate (input A, input B, output y);
    assign y = A & B;
endmodule